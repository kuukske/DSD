LIBRARY ieee;
USE ieee.std_logic_1164.all;

--///////////////////////////////////////////////////////////
--////////////////////ENTITY DECLARATION////////////////////
--/////////////////////////////////////////////////////////
ENTITY EXAMPLE_BLOCK IS

PORT
(
--CLK		:	IN	STD_LOGIC;
--NRST	:	IN	STD_LOGIC;

END EXAMPLE_BLOCK;

--///////////////////////////////////////////////////////////
--///////////////////////ARCHITECTURE///////////////////////
--/////////////////////////////////////////////////////////
ARCHITECTURE EXAMPLE_BLOCK_architecture OF EXAMPLE_BLOCK IS

BEGIN

--///////////////////////////////////////////////////////////
--//////////////////////////PROCESS/////////////////////////
--/////////////////////////////////////////////////////////
processname:	PROCESS()
	BEGIN
	END PROCESS processname;

END EXAMPLE_BLOCK_architecture;
